library verilog;
use verilog.vl_types.all;
entity tb_top_module_jpeg is
end tb_top_module_jpeg;
